
module divider_12 (

    input wire        clk,             
    input wire        rst_n,           
    input wire [10:0]  max_preset,      // ������ֵ (���ڿ��Ʒ�Ƶϵ��)


    output reg        clk_div          // ��Ƶ���ʱ�����
);

   
    reg [7:0] counter; // 8λ������

  
    always @(posedge clk or negedge rst_n) begin
        if (!rst_n) begin
            
            counter <= 8'b0;
            clk_div <= 1'b0;
        end else if (counter == max_preset) begin
            
            counter <= 8'b0;      
            clk_div <= ~clk_div;  
        end else begin
            
            counter <= counter + 1;
        end
    end

endmodule
