module tb_divider_12;

    //=========================================================================
    // 1. ��������ź�
    //=========================================================================
    reg         tb_clk;
    reg         tb_rst_n;
    reg [7:0]   tb_max_preset;

    wire        tb_clk_div;

    //=========================================================================
    // 2. ʵ��������ģ�� (DUT)
    //=========================================================================
    divider_12 u_dut (
        .clk          (tb_clk),
        .rst_n        (tb_rst_n),
        .max_preset   (tb_max_preset),
        .clk_div      (tb_clk_div)
    );

    //=========================================================================
    // 3. ����ʱ���ź� (100MHz, ����=10ns)
    //=========================================================================
    initial begin
        tb_clk = 0;
        forever #5 tb_clk = ~tb_clk;
    end

    //=========================================================================
    // 4. �������߼�
    //=========================================================================
    initial begin
        // --- ��ʼ�� ---
        tb_rst_n = 1'b0;
        tb_max_preset = 8'd0;
        $display("=================================================================");
        $display("[%0t] Testbench Started. Applying reset...", $time);
        #20;
        tb_rst_n = 1'b1; // �ͷŸ�λ
        $display("[%0t] Reset released.", $time);
        $display("=================================================================");

        // --- ���� 1: 2��Ƶ (max_preset = 0) ---
        // Ԥ��: ������� = 2 * (0+1) * 10ns = 20ns
        $display("[%0t] TEST 1: Setting max_preset = 0 (for 2x division).", $time);
        tb_max_preset = 8'd0;
        #100; // �ȴ�5���������

        // --- ���� 2: 10��Ƶ (max_preset = 4) ---
        // Ԥ��: ������� = 2 * (4+1) * 10ns = 100ns
        $display("[%0t] TEST 2: Setting max_preset = 4 (for 10x division).", $time);
        tb_max_preset = 8'd4;
        #300; // �ȴ�3���������

        // --- ���� 3: 20��Ƶ (max_preset = 9) ---
        // Ԥ��: ������� = 2 * (9+1) * 10ns = 200ns
        $display("[%0t] TEST 3: Setting max_preset = 9 (for 20x division).", $time);
        tb_max_preset = 8'd9;
        #500; // �ȴ�2.5���������

        // --- ���� 4: ��̬�л� ---
        // �Ӵ��Ƶϵ���л���С��Ƶϵ��
        $display("[%0t] TEST 4: Dynamically changing max_preset from 9 to 1.", $time);
        tb_max_preset = 8'd1; // �л���4��Ƶ
        #200; // �۲��л������Ϊ

        $display("=================================================================");
        $display("[%0t] ALL TESTS FINISHED.", $time);
        $finish;
    end

    //=========================================================================
    // 5. ������
    //=========================================================================
    // ��عؼ��źŵı仯
    initial begin
        $monitor("Time=%t | rst_n=%b | max_preset=%d | clk_div=%b", 
                 $time, tb_rst_n, tb_max_preset, tb_clk_div);
    end

endmodule