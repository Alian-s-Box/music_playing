`timescale 1ns / 1ps

//-----------------------------------------------------------------------------
// Module:      simple_button_counter_tb
// Description: simple_button_counter ģ��ļ��������ļ�
//              ���԰���������ģ3�������ܡ�
//-----------------------------------------------------------------------------
module tb_simple_button_counter;

    //=========================================================================
    // 1. ��������ź�
    //=========================================================================
    reg         tb_clk;
    reg         tb_rst_n;
    reg         tb_key_in;

    wire [1:0]  tb_count_out;

    //=========================================================================
    // 2. ʵ��������ģ�� (DUT)
    //=========================================================================
    simple_button_counter u_dut (
        .clk          (tb_clk),
        .rst_n        (tb_rst_n),
        .key_in       (tb_key_in),
        .count_out    (tb_count_out)
    );

    //=========================================================================
    // 3. ����ʱ���ź� (100MHz, ����=10ns)
    //=========================================================================
    initial begin
        tb_clk = 0;
        forever #5 tb_clk = ~tb_clk;
    end

    //=========================================================================
    // 4. ��������ģ�ⰴ������
    //=========================================================================
    // ģ��һ����Ч�İ������� (���²�����)
    task press_key;
        input integer hold_cycles; // �������ֵ�ʱ��������
        begin
            $display("[%0t] --- Simulating key press (hold for %d cycles) ---", $time, hold_cycles);
            tb_key_in = 1'b0; // �������� (�͵�ƽ)
            #(hold_cycles * 10); // ����ָ������
            tb_key_in = 1'b1; // �����ͷ� (�ߵ�ƽ)
            #100; // �ȴ�һ��ʱ����ģ�鴦��
        end
    endtask

    // ģ�ⰴ������
    task simulate_bounce;
        input integer bounce_cycles; // ������������������
        integer i;
        begin
            $display("[%0t] --- Simulating key bounce for %d ns ---", $time, bounce_cycles * 10);
            for (i = 0; i < bounce_cycles; i = i + 1) begin
                #2 tb_key_in = ~tb_key_in; // ÿ2ns��תһ�Σ�ģ���Ƶ����
            end
            tb_key_in = 1'b1; // ȷ�����������󰴼����ͷ�״̬
            #50;
        end
    endtask

    //=========================================================================
    // 5. �������߼�
    //=========================================================================
    initial begin
        // --- ��ʼ�� ---
        tb_rst_n = 1'b0;
        tb_key_in = 1'b1; // ����Ĭ��Ϊ�ߵ�ƽ��δ���£�
        $display("=================================================================");
        $display("[%0t] Testbench Started. Applying reset...", $time);
        #100;
        tb_rst_n = 1'b1; // �ͷŸ�λ
        $display("[%0t] Reset released. Initial count_out = %b", $time, tb_count_out);
        $display("=================================================================");

        // --- ���� 1: ������������֤�������� ---
        $display("[%0t] TEST 1: Normal key presses.", $time);
        press_key(200); // ����200������ (2us)��Զ��������ʱ��(160ns)
        $display("[%0t] After 1st press, count_out = %b", $time, tb_count_out);
        press_key(200);
        $display("[%0t] After 2nd press, count_out = %b", $time, tb_count_out);
        press_key(200);
        $display("[%0t] After 3rd press, count_out = %b (should be 00)", $time, tb_count_out);
        #200;

        // --- ���� 2: ������������֤�������� ---
        $display("[%0t] TEST 2: Key bounce (should be ignored).", $time);
        simulate_bounce(20); // ģ��20�ζ�������ʱ��40ns
        $display("[%0t] After bounce, count_out = %b (should be unchanged)", $time, tb_count_out);
        #200;

        // --- ���� 3: �������ȶ����£���֤���������������� ---
        $display("[%0t] TEST 3: Bounce followed by a stable press.", $time);
        simulate_bounce(20); // �ȶ���
        press_key(200);      // ���ȶ�����
        $display("[%0t] After stable press, count_out = %b (should be 01)", $time, tb_count_out);
        #200;

        // --- ���� 4: ����ʱ��̫�̣���֤�Ƿ񱻺��� ---
        $display("[%0t] TEST 4: Short key press (should be ignored).", $time);
        tb_key_in = 1'b0;
        #100; // ֻ����100ns��С����������ʱ��
        tb_key_in = 1'b1;
        $display("[%0t] After short press, count_out = %b (should be unchanged)", $time, tb_count_out);
        #200;

        $display("=================================================================");
        $display("[%0t] ALL TESTS FINISHED.", $time);
        $finish;
    end

    //=========================================================================
    // 6. ������
    //=========================================================================
    // ��عؼ��źŵı仯
    initial begin
        $monitor("Time=%t ns | rst_n=%b | key_in=%b | count_out=%b", 
                 $time, tb_rst_n, tb_key_in, tb_count_out);
    end

endmodule
