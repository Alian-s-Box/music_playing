`timescale 1ns / 1ps

//-----------------------------------------------------------------------------
// Module:      divider_clk_tb
// Description: divider_clk ģ��ļ��������ļ�
//              ��֤4��Ƶ��250,000��Ƶ���ܡ�
//-----------------------------------------------------------------------------
module tb_divider_clk;

    //=========================================================================
    // 1. ��������ź�
    //=========================================================================
    reg         tb_clk_in;
    reg         tb_rst_n;

    wire        tb_clk_div_4;
    wire        tb_clk_div_250k;

    //=========================================================================
    // 2. ʵ��������ģ�� (DUT)
    //=========================================================================
    divider_clk u_dut (
        .clk_in        (tb_clk_in),
        .rst_n         (tb_rst_n),
        .clk_div_4     (tb_clk_div_4),
        .clk_div_250k  (tb_clk_div_250k)
    );

    //=========================================================================
    // 3. ��������ʱ�� (100MHz, ����=10ns)
    //=========================================================================
    initial begin
        tb_clk_in = 0;
        forever #5 tb_clk_in = ~tb_clk_in;
    end

    //=========================================================================
    // 4. �������߼�
    //=========================================================================
    initial begin
        // --- ��ʼ�� ---
        tb_rst_n = 1'b0;
        $display("=================================================================");
        $display("[%0t] Testbench Started. Applying reset...", $time);
        #100; // ���ָ�λ100ns
        tb_rst_n = 1'b1; // �ͷŸ�λ
        $display("[%0t] Reset released.", $time);
        $display("=================================================================");

        // --- �ȴ����۲� ---
        $display("[%0t] Waiting for 3ms to observe the slow clock (clk_div_250k)...", $time);
        $display("Expected period for clk_div_4 is 40ns.");
        $display("Expected period for clk_div_250k is 2.5ms (2,500,000ns).");
        
        // �ȴ�3,000,000ns (��3ms)
        // �������� clk_div_250k ���һ���������� (2.5ms) ����ʼ��һ������
        #3_000_000;

        $display("=================================================================");
        $display("[%0t] Simulation finished. Check the waveform viewer.", $time);
        $finish;
    end

    //=========================================================================
    // 5. ������
    //=========================================================================
    // ��عؼ��źŵı仯���ر�������ʱ�ӵķ�ת
    initial begin
        $monitor("Time=%t ns | clk_div_4=%b, clk_div_250k=%b", 
                 $time, tb_clk_div_4, tb_clk_div_250k);
    end

endmodule
